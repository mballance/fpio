
`include "uvm_macros.svh"

package fpio_uvm_env_pkg;
	import uvm_pkg::*;
	import generic_sram_line_en_master_agent_pkg::*;
	import fpio_fifo_in_client_agent_pkg::*;
	import fpio_fifo_out_client_agent_pkg::*;

	`include "fpio_uvm_env.svh"
	
endpackage
