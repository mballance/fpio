
`include "uvm_macros.svh"

package fpio_env_pkg;
	import uvm_pkg::*;
	import fpio_fifo_in_client_agent_pkg::*;

	`include "fpio_env.svh"
	
endpackage
