
`include "uvm_macros.svh"

package fpio_fifo_env_pkg;
	import uvm_pkg::*;
	import fpio_fifo_in_client_agent_pkg::*;

	`include "fpio_fifo_env.svh"
	
endpackage
