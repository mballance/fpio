

`include "uvm_macros.svh"
package fpio_fifo_tests_pkg;
	import uvm_pkg::*;
	import fpio_fifo_env_pkg::*;
	
	`include "fpio_fifo_test_base.svh"
	`include "fpio_fifo_smoke_test.svh"
	
endpackage
