

`include "uvm_macros.svh"
package fpio_tests_pkg;
	import uvm_pkg::*;
	import fpio_env_pkg::*;
	
	`include "fpio_test_base.svh"
	
endpackage
